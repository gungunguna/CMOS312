*** Transient Analysis
VIN 1 0 pulse (0 5V 0ns 0ns 0ns 100ms 200ms)
R1 1 2 10K
C1 2 0 1uF
L1 2 0 1mH
.tran 0.2ms 1000ms
.control
run
plot V(1) V(2)
.endc
.end