***Pass Transistor Y = AB + C(D+E)
.subckt pass_and 1 2 3 4
M1 2 3 4 4 nmod w = 1000u l = 10u
M2 1 2 4 4 nmod w = 1000u l = 10u
.model nmod nmos level = 54 version = 4.7
.ends

.subckt pass_or 1 2 3 4
M1 2 2 4 4 nmod w = 1000u l = 10u
M2 1 3 4 4 nmod w = 1000u l = 10u
.model nmod nmos level = 54 version = 4.7
.ends

.subckt inverter 1 2 3
M1 3 1 2 2 pmod w = 1000u l = 10u
M2 3 1 0 0 nmod w = 1000u l = 10u
.model nmod nmos level = 54 version = 4.7
.model pmod pmos level = 54 version = 4.7
.ends

Va 11 0 DC 5V
Vb 12 0 DC 5V
Vc 13 0 DC 5V
Vd 14 0 DC 5V
Ve 15 0 pulse (0 5 0 0 0 10m 20m)
Vdd 2 0 DC 5V
Xb 12 2 16 inverter
Xc 13 2 20 inverter
Xe 15 2 18 inverter

Xa_and_b 11 12 16 17 pass_and
Xd_or_e 14 15 18 19 pass_or
Xdpluse_and_c 19 13 20 21 pass_and
Xdpluse_and_c_i 21 2 22 inverter
Xab_or_cdpluse 17 21 22 23 pass_or

.tran 0.1m 100m
.control
run
plot V(23) title 'Y = AB + C(D+E)' xlabel 'Time' ylabel 'Output'
.endc
.end
