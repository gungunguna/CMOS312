*** pMOS Characteristics
Vg 1 0 dc -2
Vd 3 0 dc -2.5
V1 3 2 dc 0
.model pmod pmos level = 54 version = 4.7
M1 0 1 2 2 pmod w = 100u l = 10u
.dc Vd 0 -2 -0.1
.control
run
plot i(V1) xlabel 'Vd' ylabel 'id' title 'Output char. of pMOS'
.endc
.end