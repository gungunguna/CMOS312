*** DC Analysis
VIN 1 0 5V
R1 1 2 8K
R2 2 0 2K
.dc VIN 0.0 5.0 0.1
.control
run
plot V(1) V(2)
.endc
.end