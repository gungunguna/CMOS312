*** CMOS Inverter
V1 1 0 pulse (0 5 0 0 0 10ms 20ms)
V2 2 0 DC 5V
V3 3 0 DC 0V
V4 4 0 DC 0V
Vdd 9 0 DC 5V
.model nmod nmos level = 54 version = 4.7
.model pmod pmos level = 54 version = 4.7
M1n 8 1 0 0 nmod w = 1000u l = 10u
M2n 8 2 0 0 nmod w = 1000u l = 10u
M3n 8 3 0 0 nmod w = 1000u l = 10u
M4n 8 4 0 0 nmod w = 1000u l = 10u
M1p 5 1 9 9 pmod w = 1000u l = 10u
M2p 6 2 5 5 pmod w = 1000u l = 10u
M3p 7 3 6 6 pmod w = 1000u l = 10u
M4p 8 4 7 7 pmod w = 1000u l = 10u
.tran 0.1m 100ms
.control
run
plot V(3) V(2) V(1) V(8) xlabel 'Time' ylabel 'Output' title 'CMOS Inverter'
plot V(8) xlabel 'Time' ylabel 'Output' title '4-input NOR Gate'
.endc
.end
